library verilog;
use verilog.vl_types.all;
entity Mips_tb is
end Mips_tb;
