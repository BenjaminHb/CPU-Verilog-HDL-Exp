module mips( clk, rst );

	input   clk;
	input   rst;

	wire 		RFWr;
	wire 		DMWr;
	wire 		PCWr;
	wire 		IRWr;
	wire [1:0]	EXTOp;
	wire [2:0]	ALUOp;
	wire [1:0]	NPCOp;
	wire 		BSel;
	wire 		Zero;


	assign Op =		instr[31:26];
	assign Funct =	instr[5:0];
	assign rs =		instr[25:21];
	assign rt =		instr[20:16];
	assign rd =		instr[15:11];
	assign Imm16 =	instr[15:0];
	assign IMM =	instr[25:0];


	PC U_PC (
		.clk(clk), .rst(rst), .PCWr(PCWr), .NPC(NPC), .PC(PC)
	); 

	im_4k U_IM ( 
		.addr(PC[9:0]) , .dout(im_dout)
	);


	RF U_RF (
		.A1(rs), .A2(rt), .A3(A3), .WD(WD), .clk(clk), .RFWr(RFWr), .RD1(RD1), .RD2(RD2)
	);

endmodule